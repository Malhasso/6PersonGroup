LIBRARY IEEE;
LIBRARY LPM;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE LPM.LPM_COMPONENTS.ALL;

ENTITY SRAM IS
	PORT(
		IO_CYCLE		:	IN		STD_LOGIC;
		IO_WRITE		:	IN 		STD_LOGIC;
		SRAM_ADHI_00	:	IN 		STD_LOGIC;
		SRAM_ADHI_01	:	IN 		STD_LOGIC;
		SRAM_ADHI_10	:	IN 		STD_LOGIC;
		SRAM_ADHI_11	:	IN 		STD_LOGIC;
		SRAM_DATA_EN	:	IN		STD_LOGIC;
		IO_DATA			:	INOUT	STD_LOGIC_VECTOR(15 DOWNTO 0);
		SRAM_ADDR		:	OUT		STD_LOGIC_VECTOR(17 DOWNTO 0);
		SRAM_DQ			:	INOUT	STD_LOGIC_VECTOR(15 DOWNTO 0);
		SRAM_OE_N		:	OUT		STD_LOGIC;
		SRAM_WE_N		:	OUT 	STD_LOGIC;
		SRAM_UB_N		:	OUT 	STD_LOGIC;
		SRAM_LB_N		:	OUT 	STD_LOGIC;
		SRAM_CE_N		:	OUT 	STD_LOGIC
	);
END SRAM;

ARCHITECTURE a OF SRAM IS
	TYPE STATE_TYPE IS (
		GET_ADD,
		HOLD_ADD,
		READ_SRAM,
		WRITE_SRAM,
		STANDBY
	);
	
	SIGNAL STATE		:	STATE_TYPE;
	SIGNAL IO_READ		:	STD_LOGIC;
	SIGNAL FULL_ADDR	:	STD_LOGIC_VECTOR(17 DOWNTO 0);
	SIGNAL SRAM_EN		:	STD_LOGIC;
	SIGNAL ADDR_EN		:	STD_LOGIC;
	SIGNAL ADDRESS_LOW	:	STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL ADDRESS_HI	:	STD_LOGIC_VECTOR(1 DOWNTO 0);
	SIGNAL SRAM_CTRL	:	STD_LOGIC_VECTOR(1 DOWNTO 0);


BEGIN
	IO_BUS: lpm_bustri
	GENERIC MAP (
		lpm_width => 16
	)
	PORT MAP (
	data 	 	=> 	IO_DATA,
	enabledt	=>	IO_WRITE,
	tridata 	=>	SRAM_DQ,
	enabletr	=>	IO_READ,
	result		=>	IO_DATA
	);
	
	IO_READ 	<= (NOT(IO_WRITE) AND IO_CYCLE);
	
	PROCESS(IO_WRITE, IO_CYCLE)
	BEGIN
		IF (SRAM_EN = '0') THEN
			STATE <= STANDBY;
		ELSIF (SRAM_EN = '1') THEN
			CASE STATE IS
				WHEN STANDBY =>
					IF (ADDR_EN = '1') THEN
						STATE <= GET_ADD;
					ELSIF (SRAM_DATA_EN = '1') THEN
						IF ( IO_READ = '1') THEN
							STATE <= READ_SRAM;
						ELSIF ( IO_WRITE = '1') THEN
							STATE <= WRITE_SRAM;
						END IF;
					ELSE
						STATE <= STANDBY;
					END IF;
				WHEN GET_ADD =>
					IF ((SRAM_ADHI_00 = '1') AND (IO_CYCLE = '1') AND (IO_WRITE = '1')) THEN
						FULL_ADDR <= "00" & IO_DATA;
						STATE <= HOLD_ADD;
					ELSIF ((SRAM_ADHI_01 = '1') AND (IO_CYCLE = '1') AND (IO_WRITE = '1')) THEN
						FULL_ADDR <= "01" & IO_DATA;
						STATE <= HOLD_ADD;
					ELSIF ((SRAM_ADHI_10 = '1') AND (IO_CYCLE = '1') AND (IO_WRITE = '1')) THEN
						FULL_ADDR <= "10" & IO_DATA;
						STATE <= HOLD_ADD;
					ELSIF ((SRAM_ADHI_11 = '1') AND (IO_CYCLE = '1') AND (IO_WRITE = '1')) THEN
						FULL_ADDR <= "11" & IO_DATA;
						STATE <= HOLD_ADD;
					ELSE
						STATE <= GET_ADD;
					END IF;
				WHEN READ_SRAM =>
					STATE <= STANDBY;
				WHEN WRITE_SRAM =>
					STATE <= STANDBY;
				WHEN HOLD_ADD =>
					IF (ADDR_EN = '1') THEN
						STATE <= HOLD_ADD;
					ELSE
						STATE <= STANDBY;
					END IF;
				WHEN OTHERS =>
					STATE <= STANDBY;
			END CASE;	
		END IF;
	END PROCESS;
	
	WITH STATE SELECT
		SRAM_OE_N <= '0' WHEN READ_SRAM,
					 '1' WHEN OTHERS;
	WITH STATE SELECT
		SRAM_WE_N <= '0' WHEN WRITE_SRAM,
					 '1' WHEN OTHERS;
	
	SRAM_ADDR <= FULL_ADDR;
				  
	SRAM_UB_N <= '0';
	SRAM_LB_N <= '0';
	SRAM_CE_N <= '0';
			
	SRAM_EN		<= (IO_WRITE OR IO_CYCLE);
	ADDR_EN		<= (SRAM_ADHI_00  OR SRAM_ADHI_01 OR SRAM_ADHI_10 OR SRAM_ADHI_11);
END a;	




	